library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.all;

entity registros is
    Port ( CLK : in  STD_LOGIC;
           WE3 : in  STD_LOGIC; -- ENABLER
           A1 : in  STD_LOGIC_VECTOR (4 downto 0);
           A2 : in  STD_LOGIC_VECTOR (4 downto 0);
           A3 : in  STD_LOGIC_VECTOR (4 downto 0);
           WD3 : in  STD_LOGIC_VECTOR (31 downto 0);	-- DATO A ESCRIBIR
           RD1 : out  STD_LOGIC_VECTOR (31 downto 0);
           RD2 : out  STD_LOGIC_VECTOR (31 downto 0));
end registros;

architecture arch_registros of registros is
type ramtype is array (0 to 31) of STD_LOGIC_VECTOR(31 downto 0);
signal mem: ramtype:= (
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000000000",
	"00000000000000000000000000101110", ---$29 Stack Pointer (46) deja 2 lugares de 32 bits: 1 para el controlador de boton y 1 para LCD
	"00000000000000000000000000000000",
	"00000000000000000000000000000000"--ra
	--OTHERS => "00000000000000000000000000000000"
);

begin
	-- ESPERAMOS EL CLOCK
	process(CLK,WD3,A3,A2,A1,mem)	-- PROCESO PARA ESCRIBIR EL DATO EN LA DIRECCION A3
	begin
		if (CLK'event and CLK = '1' and WE3 = '1' ) then
			mem(conv_integer(A3)) <= WD3;
		end if;
	 
	
	if(conv_integer(A1) = 0) then
		RD1 <= X"00000000"; --EL REGISTRO 0 SIEMPRE TIENE 0 ADENTRO
	else
		RD1 <= mem(conv_integer(A1)); -- SI NO ES CERO PONGO EL DATO
	end if;
	if(conv_integer(A2) = 0) then -- HACES LO MISMO PARA A2
		RD2 <= X"00000000";
	else
		RD2 <= mem(conv_integer(A2));
	end if;
	end process;
end arch_registros;

